/*
-Practico 1
-Ejercicio 6

Decodificador para generar las seniales de control

*/
`include "macros.sv"

module maindec (
    input  logic [10:0] Op,
    output logic        Reg2Loc,
    output logic        ALUSrc,
    output logic        MemtoReg,
    output logic        RegWrite,
    output logic        MemRead,
    output logic        MemWrite,
    output logic        Branch,
    output logic [1:0]  ALUOp,
    output logic        Uncondbranch,
    output logic        BranchSrc
);

    always_comb
    begin
        Uncondbranch = 1'b0;
        BranchSrc    = 1'b0;

        casez(Op)
            `LDUR: begin
                Reg2Loc  = 1'b0;
                ALUSrc   = 1'b1;
                MemtoReg = 1'b1;
                RegWrite = 1'b1;
                MemRead  = 1'b1;
                MemWrite = 1'b0;
                Branch   = 1'b0;
                ALUOp    = 2'b00;
            end

            `STUR: begin
                Reg2Loc  = 1'b1;
                ALUSrc   = 1'b1;
                MemtoReg = 1'b0;
                RegWrite = 1'b0;
                MemRead  = 1'b0;
                MemWrite = 1'b1;
                Branch   = 1'b0;
                ALUOp    = 2'b00;
            end

            `CBZ: begin
                Reg2Loc  = 1'b1;
                ALUSrc   = 1'b0;
                MemtoReg = 1'b0;
                RegWrite = 1'b0;
                MemRead  = 1'b0;
                MemWrite = 1'b0;
                Branch   = 1'b1;
                ALUOp    = 2'b01;
            end

            `ADD: begin
                Reg2Loc  = 1'b0;
                ALUSrc   = 1'b0;
                MemtoReg = 1'b0;
                RegWrite = 1'b1;
                MemRead  = 1'b0;
                MemWrite = 1'b0;
                Branch   = 1'b0;
                ALUOp    = 2'b10;
            end

            `SUB: begin
                Reg2Loc  = 1'b0;
                ALUSrc   = 1'b0;
                MemtoReg = 1'b0;
                RegWrite = 1'b1;
                MemRead  = 1'b0;
                MemWrite = 1'b0;
                Branch   = 1'b0;
                ALUOp    = 2'b10;
            end

            `AND: begin
                Reg2Loc  = 1'b0;
                ALUSrc   = 1'b0;
                MemtoReg = 1'b0;
                RegWrite = 1'b1;
                MemRead  = 1'b0;
                MemWrite = 1'b0;
                Branch   = 1'b0;
                ALUOp    = 2'b10;
            end

            `ORR: begin
                Reg2Loc  = 1'b0;
                ALUSrc   = 1'b0;
                MemtoReg = 1'b0;
                RegWrite = 1'b1;
                MemRead  = 1'b0;
                MemWrite = 1'b0;
                Branch   = 1'b0;
                ALUOp    = 2'b10;
            end

            `B: begin
                Reg2Loc      = 1'b0;
                ALUSrc       = 1'b0;
                MemtoReg     = 1'b0;
                RegWrite     = 1'b0;
                MemRead      = 1'b0;
                MemWrite     = 1'b0;
                Branch       = 1'b0;
                ALUOp        = 2'b00;
                Uncondbranch = 1'b1;
            end

            `BR: begin
                Reg2Loc      = 1'b0;
                ALUSrc       = 1'b0;
                MemtoReg     = 1'b0;
                RegWrite     = 1'b0;
                MemRead      = 1'b0;
                MemWrite     = 1'b0;
                Branch       = 1'b0;
                ALUOp        = 2'b00;
                Uncondbranch = 1'b1;
                BranchSrc    = 1'b1;
            end

            default: begin           // undefined opcode (all at 0)
                Reg2Loc  = 1'b0;
                ALUSrc   = 1'b0;
                MemtoReg = 1'b0;
                RegWrite = 1'b0;
                MemRead  = 1'b0;
                MemWrite = 1'b0;
                Branch   = 1'b0;
                ALUOp    = 2'b00;
            end
        endcase
    end

endmodule
